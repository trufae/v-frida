module host

#flag -Iext/frida
#flag -Lext/frida
#flag -lfrida-core -lresolv -framework Foundation -lbsm -framework AppKit

#include <frida-core.h>


