module host

#flag -Iext/frida
#flag ext/frida/libfrida-core.a -lresolv -framework Foundation -lbsm -framework AppKit

#include <frida-core.h>


