module frida
